
module eindopdracht (
	clk_clk,
	pio_buttons_external_connection_export,
	pio_switches_external_connection_export,
	rgb_framebuffer_0_rgb_matrix_conduit_r1,
	rgb_framebuffer_0_rgb_matrix_conduit_g1,
	rgb_framebuffer_0_rgb_matrix_conduit_b1,
	rgb_framebuffer_0_rgb_matrix_conduit_r2,
	rgb_framebuffer_0_rgb_matrix_conduit_g2,
	rgb_framebuffer_0_rgb_matrix_conduit_b2,
	rgb_framebuffer_0_rgb_matrix_conduit_addr_a,
	rgb_framebuffer_0_rgb_matrix_conduit_addr_b,
	rgb_framebuffer_0_rgb_matrix_conduit_addr_c,
	rgb_framebuffer_0_rgb_matrix_conduit_clk_out,
	rgb_framebuffer_0_rgb_matrix_conduit_lat,
	rgb_framebuffer_0_rgb_matrix_conduit_oe_n);	

	input		clk_clk;
	input	[3:0]	pio_buttons_external_connection_export;
	input	[9:0]	pio_switches_external_connection_export;
	output		rgb_framebuffer_0_rgb_matrix_conduit_r1;
	output		rgb_framebuffer_0_rgb_matrix_conduit_g1;
	output		rgb_framebuffer_0_rgb_matrix_conduit_b1;
	output		rgb_framebuffer_0_rgb_matrix_conduit_r2;
	output		rgb_framebuffer_0_rgb_matrix_conduit_g2;
	output		rgb_framebuffer_0_rgb_matrix_conduit_b2;
	output		rgb_framebuffer_0_rgb_matrix_conduit_addr_a;
	output		rgb_framebuffer_0_rgb_matrix_conduit_addr_b;
	output		rgb_framebuffer_0_rgb_matrix_conduit_addr_c;
	output		rgb_framebuffer_0_rgb_matrix_conduit_clk_out;
	output		rgb_framebuffer_0_rgb_matrix_conduit_lat;
	output		rgb_framebuffer_0_rgb_matrix_conduit_oe_n;
endmodule
