-- eindopdracht.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity eindopdracht is
	port (
		clk_clk                : in  std_logic                     := '0';             --           clk.clk
		matrix_output_readdata : out std_logic_vector(31 downto 0);                    -- matrix_output.readdata
		pio_buttons_export     : in  std_logic_vector(3 downto 0)  := (others => '0'); --   pio_buttons.export
		pio_leds_export        : out std_logic_vector(9 downto 0);                     --      pio_leds.export
		pio_switches_export    : in  std_logic_vector(9 downto 0)  := (others => '0')  --  pio_switches.export
	);
end entity eindopdracht;

architecture rtl of eindopdracht is
	component eindopdracht_JTAG_DEBUG is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component eindopdracht_JTAG_DEBUG;

	component eindopdracht_Processor_Nios is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(19 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(19 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component eindopdracht_Processor_Nios;

	component eindopdracht_RAM is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component eindopdracht_RAM;

	component reg32_avalon_interface is
		port (
			reset      : in  std_logic                     := 'X';             -- reset
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			Q_export   : out std_logic_vector(31 downto 0);                    -- readdata
			clock      : in  std_logic                     := 'X'              -- clk
		);
	end component reg32_avalon_interface;

	component eindopdracht_performance_checker_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component eindopdracht_performance_checker_0;

	component eindopdracht_pio_buttons is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component eindopdracht_pio_buttons;

	component eindopdracht_pio_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component eindopdracht_pio_leds;

	component eindopdracht_pio_switches is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component eindopdracht_pio_switches;

	component eindopdracht_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component eindopdracht_sysid_qsys_0;

	component eindopdracht_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component eindopdracht_timer_0;

	component eindopdracht_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                      : in  std_logic                     := 'X';             -- clk
			Processor_Nios_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Processor_Nios_data_master_address                 : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			Processor_Nios_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			Processor_Nios_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			Processor_Nios_data_master_read                    : in  std_logic                     := 'X';             -- read
			Processor_Nios_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			Processor_Nios_data_master_write                   : in  std_logic                     := 'X';             -- write
			Processor_Nios_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Processor_Nios_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			Processor_Nios_instruction_master_address          : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			Processor_Nios_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			Processor_Nios_instruction_master_read             : in  std_logic                     := 'X';             -- read
			Processor_Nios_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			JTAG_DEBUG_avalon_jtag_slave_address               : out std_logic_vector(0 downto 0);                     -- address
			JTAG_DEBUG_avalon_jtag_slave_write                 : out std_logic;                                        -- write
			JTAG_DEBUG_avalon_jtag_slave_read                  : out std_logic;                                        -- read
			JTAG_DEBUG_avalon_jtag_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_DEBUG_avalon_jtag_slave_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_DEBUG_avalon_jtag_slave_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			JTAG_DEBUG_avalon_jtag_slave_chipselect            : out std_logic;                                        -- chipselect
			led_matrix_0_avalon_slave_0_address                : out std_logic_vector(1 downto 0);                     -- address
			led_matrix_0_avalon_slave_0_write                  : out std_logic;                                        -- write
			led_matrix_0_avalon_slave_0_read                   : out std_logic;                                        -- read
			led_matrix_0_avalon_slave_0_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_matrix_0_avalon_slave_0_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			led_matrix_0_avalon_slave_0_byteenable             : out std_logic_vector(3 downto 0);                     -- byteenable
			led_matrix_0_avalon_slave_0_chipselect             : out std_logic;                                        -- chipselect
			performance_checker_0_control_slave_address        : out std_logic_vector(3 downto 0);                     -- address
			performance_checker_0_control_slave_write          : out std_logic;                                        -- write
			performance_checker_0_control_slave_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			performance_checker_0_control_slave_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			performance_checker_0_control_slave_begintransfer  : out std_logic;                                        -- begintransfer
			pio_buttons_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			pio_buttons_s1_write                               : out std_logic;                                        -- write
			pio_buttons_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_buttons_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			pio_buttons_s1_chipselect                          : out std_logic;                                        -- chipselect
			pio_leds_s1_address                                : out std_logic_vector(1 downto 0);                     -- address
			pio_leds_s1_write                                  : out std_logic;                                        -- write
			pio_leds_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_leds_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			pio_leds_s1_chipselect                             : out std_logic;                                        -- chipselect
			pio_switches_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			pio_switches_s1_write                              : out std_logic;                                        -- write
			pio_switches_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_switches_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			pio_switches_s1_chipselect                         : out std_logic;                                        -- chipselect
			Processor_Nios_jtag_debug_module_address           : out std_logic_vector(8 downto 0);                     -- address
			Processor_Nios_jtag_debug_module_write             : out std_logic;                                        -- write
			Processor_Nios_jtag_debug_module_read              : out std_logic;                                        -- read
			Processor_Nios_jtag_debug_module_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Processor_Nios_jtag_debug_module_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			Processor_Nios_jtag_debug_module_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			Processor_Nios_jtag_debug_module_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			Processor_Nios_jtag_debug_module_debugaccess       : out std_logic;                                        -- debugaccess
			RAM_s1_address                                     : out std_logic_vector(15 downto 0);                    -- address
			RAM_s1_write                                       : out std_logic;                                        -- write
			RAM_s1_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			RAM_s1_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			RAM_s1_byteenable                                  : out std_logic_vector(3 downto 0);                     -- byteenable
			RAM_s1_chipselect                                  : out std_logic;                                        -- chipselect
			RAM_s1_clken                                       : out std_logic;                                        -- clken
			sysid_qsys_0_control_slave_address                 : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                                 : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                   : out std_logic;                                        -- write
			timer_0_s1_readdata                                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                               : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                              : out std_logic                                         -- chipselect
		);
	end component eindopdracht_mm_interconnect_0;

	component eindopdracht_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component eindopdracht_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal processor_nios_jtag_debug_module_reset_reset                        : std_logic;                     -- Processor_Nios:jtag_debug_module_resetrequest -> rst_controller:reset_in0
	signal processor_nios_data_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor_Nios_data_master_readdata -> Processor_Nios:d_readdata
	signal processor_nios_data_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:Processor_Nios_data_master_waitrequest -> Processor_Nios:d_waitrequest
	signal processor_nios_data_master_debugaccess                              : std_logic;                     -- Processor_Nios:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:Processor_Nios_data_master_debugaccess
	signal processor_nios_data_master_address                                  : std_logic_vector(19 downto 0); -- Processor_Nios:d_address -> mm_interconnect_0:Processor_Nios_data_master_address
	signal processor_nios_data_master_byteenable                               : std_logic_vector(3 downto 0);  -- Processor_Nios:d_byteenable -> mm_interconnect_0:Processor_Nios_data_master_byteenable
	signal processor_nios_data_master_read                                     : std_logic;                     -- Processor_Nios:d_read -> mm_interconnect_0:Processor_Nios_data_master_read
	signal processor_nios_data_master_write                                    : std_logic;                     -- Processor_Nios:d_write -> mm_interconnect_0:Processor_Nios_data_master_write
	signal processor_nios_data_master_writedata                                : std_logic_vector(31 downto 0); -- Processor_Nios:d_writedata -> mm_interconnect_0:Processor_Nios_data_master_writedata
	signal processor_nios_instruction_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor_Nios_instruction_master_readdata -> Processor_Nios:i_readdata
	signal processor_nios_instruction_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:Processor_Nios_instruction_master_waitrequest -> Processor_Nios:i_waitrequest
	signal processor_nios_instruction_master_address                           : std_logic_vector(19 downto 0); -- Processor_Nios:i_address -> mm_interconnect_0:Processor_Nios_instruction_master_address
	signal processor_nios_instruction_master_read                              : std_logic;                     -- Processor_Nios:i_read -> mm_interconnect_0:Processor_Nios_instruction_master_read
	signal mm_interconnect_0_jtag_debug_avalon_jtag_slave_chipselect           : std_logic;                     -- mm_interconnect_0:JTAG_DEBUG_avalon_jtag_slave_chipselect -> JTAG_DEBUG:av_chipselect
	signal mm_interconnect_0_jtag_debug_avalon_jtag_slave_readdata             : std_logic_vector(31 downto 0); -- JTAG_DEBUG:av_readdata -> mm_interconnect_0:JTAG_DEBUG_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_debug_avalon_jtag_slave_waitrequest          : std_logic;                     -- JTAG_DEBUG:av_waitrequest -> mm_interconnect_0:JTAG_DEBUG_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_debug_avalon_jtag_slave_address              : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_DEBUG_avalon_jtag_slave_address -> JTAG_DEBUG:av_address
	signal mm_interconnect_0_jtag_debug_avalon_jtag_slave_read                 : std_logic;                     -- mm_interconnect_0:JTAG_DEBUG_avalon_jtag_slave_read -> mm_interconnect_0_jtag_debug_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_debug_avalon_jtag_slave_write                : std_logic;                     -- mm_interconnect_0:JTAG_DEBUG_avalon_jtag_slave_write -> mm_interconnect_0_jtag_debug_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_debug_avalon_jtag_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_DEBUG_avalon_jtag_slave_writedata -> JTAG_DEBUG:av_writedata
	signal mm_interconnect_0_led_matrix_0_avalon_slave_0_chipselect            : std_logic;                     -- mm_interconnect_0:led_matrix_0_avalon_slave_0_chipselect -> led_matrix_0:chipselect
	signal mm_interconnect_0_led_matrix_0_avalon_slave_0_readdata              : std_logic_vector(31 downto 0); -- led_matrix_0:readdata -> mm_interconnect_0:led_matrix_0_avalon_slave_0_readdata
	signal mm_interconnect_0_led_matrix_0_avalon_slave_0_address               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_matrix_0_avalon_slave_0_address -> led_matrix_0:address
	signal mm_interconnect_0_led_matrix_0_avalon_slave_0_read                  : std_logic;                     -- mm_interconnect_0:led_matrix_0_avalon_slave_0_read -> led_matrix_0:read
	signal mm_interconnect_0_led_matrix_0_avalon_slave_0_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:led_matrix_0_avalon_slave_0_byteenable -> led_matrix_0:byteenable
	signal mm_interconnect_0_led_matrix_0_avalon_slave_0_write                 : std_logic;                     -- mm_interconnect_0:led_matrix_0_avalon_slave_0_write -> led_matrix_0:write
	signal mm_interconnect_0_led_matrix_0_avalon_slave_0_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_matrix_0_avalon_slave_0_writedata -> led_matrix_0:writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata               : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_performance_checker_0_control_slave_readdata      : std_logic_vector(31 downto 0); -- performance_checker_0:readdata -> mm_interconnect_0:performance_checker_0_control_slave_readdata
	signal mm_interconnect_0_performance_checker_0_control_slave_address       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:performance_checker_0_control_slave_address -> performance_checker_0:address
	signal mm_interconnect_0_performance_checker_0_control_slave_begintransfer : std_logic;                     -- mm_interconnect_0:performance_checker_0_control_slave_begintransfer -> performance_checker_0:begintransfer
	signal mm_interconnect_0_performance_checker_0_control_slave_write         : std_logic;                     -- mm_interconnect_0:performance_checker_0_control_slave_write -> performance_checker_0:write
	signal mm_interconnect_0_performance_checker_0_control_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:performance_checker_0_control_slave_writedata -> performance_checker_0:writedata
	signal mm_interconnect_0_processor_nios_jtag_debug_module_readdata         : std_logic_vector(31 downto 0); -- Processor_Nios:jtag_debug_module_readdata -> mm_interconnect_0:Processor_Nios_jtag_debug_module_readdata
	signal mm_interconnect_0_processor_nios_jtag_debug_module_waitrequest      : std_logic;                     -- Processor_Nios:jtag_debug_module_waitrequest -> mm_interconnect_0:Processor_Nios_jtag_debug_module_waitrequest
	signal mm_interconnect_0_processor_nios_jtag_debug_module_debugaccess      : std_logic;                     -- mm_interconnect_0:Processor_Nios_jtag_debug_module_debugaccess -> Processor_Nios:jtag_debug_module_debugaccess
	signal mm_interconnect_0_processor_nios_jtag_debug_module_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:Processor_Nios_jtag_debug_module_address -> Processor_Nios:jtag_debug_module_address
	signal mm_interconnect_0_processor_nios_jtag_debug_module_read             : std_logic;                     -- mm_interconnect_0:Processor_Nios_jtag_debug_module_read -> Processor_Nios:jtag_debug_module_read
	signal mm_interconnect_0_processor_nios_jtag_debug_module_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Processor_Nios_jtag_debug_module_byteenable -> Processor_Nios:jtag_debug_module_byteenable
	signal mm_interconnect_0_processor_nios_jtag_debug_module_write            : std_logic;                     -- mm_interconnect_0:Processor_Nios_jtag_debug_module_write -> Processor_Nios:jtag_debug_module_write
	signal mm_interconnect_0_processor_nios_jtag_debug_module_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Processor_Nios_jtag_debug_module_writedata -> Processor_Nios:jtag_debug_module_writedata
	signal mm_interconnect_0_ram_s1_chipselect                                 : std_logic;                     -- mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	signal mm_interconnect_0_ram_s1_readdata                                   : std_logic_vector(31 downto 0); -- RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	signal mm_interconnect_0_ram_s1_address                                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:RAM_s1_address -> RAM:address
	signal mm_interconnect_0_ram_s1_byteenable                                 : std_logic_vector(3 downto 0);  -- mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	signal mm_interconnect_0_ram_s1_write                                      : std_logic;                     -- mm_interconnect_0:RAM_s1_write -> RAM:write
	signal mm_interconnect_0_ram_s1_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	signal mm_interconnect_0_ram_s1_clken                                      : std_logic;                     -- mm_interconnect_0:RAM_s1_clken -> RAM:clken
	signal mm_interconnect_0_pio_buttons_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:pio_buttons_s1_chipselect -> pio_buttons:chipselect
	signal mm_interconnect_0_pio_buttons_s1_readdata                           : std_logic_vector(31 downto 0); -- pio_buttons:readdata -> mm_interconnect_0:pio_buttons_s1_readdata
	signal mm_interconnect_0_pio_buttons_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_buttons_s1_address -> pio_buttons:address
	signal mm_interconnect_0_pio_buttons_s1_write                              : std_logic;                     -- mm_interconnect_0:pio_buttons_s1_write -> mm_interconnect_0_pio_buttons_s1_write:in
	signal mm_interconnect_0_pio_buttons_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_buttons_s1_writedata -> pio_buttons:writedata
	signal mm_interconnect_0_pio_switches_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:pio_switches_s1_chipselect -> pio_switches:chipselect
	signal mm_interconnect_0_pio_switches_s1_readdata                          : std_logic_vector(31 downto 0); -- pio_switches:readdata -> mm_interconnect_0:pio_switches_s1_readdata
	signal mm_interconnect_0_pio_switches_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_switches_s1_address -> pio_switches:address
	signal mm_interconnect_0_pio_switches_s1_write                             : std_logic;                     -- mm_interconnect_0:pio_switches_s1_write -> mm_interconnect_0_pio_switches_s1_write:in
	signal mm_interconnect_0_pio_switches_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_switches_s1_writedata -> pio_switches:writedata
	signal mm_interconnect_0_timer_0_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                               : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                                : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                                  : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                              : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_pio_leds_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:pio_leds_s1_chipselect -> pio_leds:chipselect
	signal mm_interconnect_0_pio_leds_s1_readdata                              : std_logic_vector(31 downto 0); -- pio_leds:readdata -> mm_interconnect_0:pio_leds_s1_readdata
	signal mm_interconnect_0_pio_leds_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_leds_s1_address -> pio_leds:address
	signal mm_interconnect_0_pio_leds_s1_write                                 : std_logic;                     -- mm_interconnect_0:pio_leds_s1_write -> mm_interconnect_0_pio_leds_s1_write:in
	signal mm_interconnect_0_pio_leds_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_leds_s1_writedata -> pio_leds:writedata
	signal irq_mapper_receiver0_irq                                            : std_logic;                     -- JTAG_DEBUG:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                            : std_logic;                     -- timer_0:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                            : std_logic;                     -- pio_buttons:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                            : std_logic;                     -- pio_switches:irq -> irq_mapper:receiver3_irq
	signal processor_nios_d_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> Processor_Nios:d_irq
	signal rst_controller_reset_out_reset                                      : std_logic;                     -- rst_controller:reset_out -> [RAM:reset, irq_mapper:reset, led_matrix_0:reset, mm_interconnect_0:Processor_Nios_reset_n_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                  : std_logic;                     -- rst_controller:reset_req -> [Processor_Nios:reset_req, RAM:reset_req, rst_translator:reset_req_in]
	signal mm_interconnect_0_jtag_debug_avalon_jtag_slave_read_ports_inv       : std_logic;                     -- mm_interconnect_0_jtag_debug_avalon_jtag_slave_read:inv -> JTAG_DEBUG:av_read_n
	signal mm_interconnect_0_jtag_debug_avalon_jtag_slave_write_ports_inv      : std_logic;                     -- mm_interconnect_0_jtag_debug_avalon_jtag_slave_write:inv -> JTAG_DEBUG:av_write_n
	signal mm_interconnect_0_pio_buttons_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_pio_buttons_s1_write:inv -> pio_buttons:write_n
	signal mm_interconnect_0_pio_switches_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_pio_switches_s1_write:inv -> pio_switches:write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_pio_leds_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_pio_leds_s1_write:inv -> pio_leds:write_n
	signal rst_controller_reset_out_reset_ports_inv                            : std_logic;                     -- rst_controller_reset_out_reset:inv -> [JTAG_DEBUG:rst_n, Processor_Nios:reset_n, performance_checker_0:reset_n, pio_buttons:reset_n, pio_leds:reset_n, pio_switches:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n]

begin

	jtag_debug : component eindopdracht_JTAG_DEBUG
		port map (
			clk            => clk_clk,                                                        --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                       --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_debug_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_debug_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_debug_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_debug_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_debug_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_debug_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_debug_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                        --               irq.irq
		);

	processor_nios : component eindopdracht_Processor_Nios
		port map (
			clk                                   => clk_clk,                                                        --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                       --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                             --                          .reset_req
			d_address                             => processor_nios_data_master_address,                             --               data_master.address
			d_byteenable                          => processor_nios_data_master_byteenable,                          --                          .byteenable
			d_read                                => processor_nios_data_master_read,                                --                          .read
			d_readdata                            => processor_nios_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => processor_nios_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => processor_nios_data_master_write,                               --                          .write
			d_writedata                           => processor_nios_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => processor_nios_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => processor_nios_instruction_master_address,                      --        instruction_master.address
			i_read                                => processor_nios_instruction_master_read,                         --                          .read
			i_readdata                            => processor_nios_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => processor_nios_instruction_master_waitrequest,                  --                          .waitrequest
			d_irq                                 => processor_nios_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => processor_nios_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_processor_nios_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_processor_nios_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_processor_nios_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_processor_nios_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_processor_nios_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_processor_nios_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_processor_nios_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_processor_nios_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                            -- custom_instruction_master.readra
		);

	ram : component eindopdracht_RAM
		port map (
			clk        => clk_clk,                             --   clk1.clk
			address    => mm_interconnect_0_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,      -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,  --       .reset_req
			freeze     => '0'                                  -- (terminated)
		);

	led_matrix_0 : component reg32_avalon_interface
		port map (
			reset      => rst_controller_reset_out_reset,                           --    clock_reset.reset
			read       => mm_interconnect_0_led_matrix_0_avalon_slave_0_read,       -- avalon_slave_0.read
			write      => mm_interconnect_0_led_matrix_0_avalon_slave_0_write,      --               .write
			chipselect => mm_interconnect_0_led_matrix_0_avalon_slave_0_chipselect, --               .chipselect
			readdata   => mm_interconnect_0_led_matrix_0_avalon_slave_0_readdata,   --               .readdata
			writedata  => mm_interconnect_0_led_matrix_0_avalon_slave_0_writedata,  --               .writedata
			byteenable => mm_interconnect_0_led_matrix_0_avalon_slave_0_byteenable, --               .byteenable
			address    => mm_interconnect_0_led_matrix_0_avalon_slave_0_address,    --               .address
			Q_export   => matrix_output_readdata,                                   --    conduit_end.readdata
			clock      => clk_clk                                                   --     clock_sink.clk
		);

	performance_checker_0 : component eindopdracht_performance_checker_0
		port map (
			clk           => clk_clk,                                                             --           clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                            --         reset.reset_n
			address       => mm_interconnect_0_performance_checker_0_control_slave_address,       -- control_slave.address
			begintransfer => mm_interconnect_0_performance_checker_0_control_slave_begintransfer, --              .begintransfer
			readdata      => mm_interconnect_0_performance_checker_0_control_slave_readdata,      --              .readdata
			write         => mm_interconnect_0_performance_checker_0_control_slave_write,         --              .write
			writedata     => mm_interconnect_0_performance_checker_0_control_slave_writedata      --              .writedata
		);

	pio_buttons : component eindopdracht_pio_buttons
		port map (
			clk        => clk_clk,                                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_pio_buttons_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_buttons_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_buttons_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_buttons_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_buttons_s1_readdata,        --                    .readdata
			in_port    => pio_buttons_export,                               -- external_connection.export
			irq        => irq_mapper_receiver2_irq                          --                 irq.irq
		);

	pio_leds : component eindopdracht_pio_leds
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_pio_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_leds_s1_readdata,        --                    .readdata
			out_port   => pio_leds_export                                -- external_connection.export
		);

	pio_switches : component eindopdracht_pio_switches
		port map (
			clk        => clk_clk,                                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_pio_switches_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_switches_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_switches_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_switches_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_switches_s1_readdata,        --                    .readdata
			in_port    => pio_switches_export,                               -- external_connection.export
			irq        => irq_mapper_receiver3_irq                           --                 irq.irq
		);

	sysid_qsys_0 : component eindopdracht_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	timer_0 : component eindopdracht_timer_0
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                      --   irq.irq
		);

	mm_interconnect_0 : component eindopdracht_mm_interconnect_0
		port map (
			clk_0_clk_clk                                      => clk_clk,                                                             --                                    clk_0_clk.clk
			Processor_Nios_reset_n_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                      -- Processor_Nios_reset_n_reset_bridge_in_reset.reset
			Processor_Nios_data_master_address                 => processor_nios_data_master_address,                                  --                   Processor_Nios_data_master.address
			Processor_Nios_data_master_waitrequest             => processor_nios_data_master_waitrequest,                              --                                             .waitrequest
			Processor_Nios_data_master_byteenable              => processor_nios_data_master_byteenable,                               --                                             .byteenable
			Processor_Nios_data_master_read                    => processor_nios_data_master_read,                                     --                                             .read
			Processor_Nios_data_master_readdata                => processor_nios_data_master_readdata,                                 --                                             .readdata
			Processor_Nios_data_master_write                   => processor_nios_data_master_write,                                    --                                             .write
			Processor_Nios_data_master_writedata               => processor_nios_data_master_writedata,                                --                                             .writedata
			Processor_Nios_data_master_debugaccess             => processor_nios_data_master_debugaccess,                              --                                             .debugaccess
			Processor_Nios_instruction_master_address          => processor_nios_instruction_master_address,                           --            Processor_Nios_instruction_master.address
			Processor_Nios_instruction_master_waitrequest      => processor_nios_instruction_master_waitrequest,                       --                                             .waitrequest
			Processor_Nios_instruction_master_read             => processor_nios_instruction_master_read,                              --                                             .read
			Processor_Nios_instruction_master_readdata         => processor_nios_instruction_master_readdata,                          --                                             .readdata
			JTAG_DEBUG_avalon_jtag_slave_address               => mm_interconnect_0_jtag_debug_avalon_jtag_slave_address,              --                 JTAG_DEBUG_avalon_jtag_slave.address
			JTAG_DEBUG_avalon_jtag_slave_write                 => mm_interconnect_0_jtag_debug_avalon_jtag_slave_write,                --                                             .write
			JTAG_DEBUG_avalon_jtag_slave_read                  => mm_interconnect_0_jtag_debug_avalon_jtag_slave_read,                 --                                             .read
			JTAG_DEBUG_avalon_jtag_slave_readdata              => mm_interconnect_0_jtag_debug_avalon_jtag_slave_readdata,             --                                             .readdata
			JTAG_DEBUG_avalon_jtag_slave_writedata             => mm_interconnect_0_jtag_debug_avalon_jtag_slave_writedata,            --                                             .writedata
			JTAG_DEBUG_avalon_jtag_slave_waitrequest           => mm_interconnect_0_jtag_debug_avalon_jtag_slave_waitrequest,          --                                             .waitrequest
			JTAG_DEBUG_avalon_jtag_slave_chipselect            => mm_interconnect_0_jtag_debug_avalon_jtag_slave_chipselect,           --                                             .chipselect
			led_matrix_0_avalon_slave_0_address                => mm_interconnect_0_led_matrix_0_avalon_slave_0_address,               --                  led_matrix_0_avalon_slave_0.address
			led_matrix_0_avalon_slave_0_write                  => mm_interconnect_0_led_matrix_0_avalon_slave_0_write,                 --                                             .write
			led_matrix_0_avalon_slave_0_read                   => mm_interconnect_0_led_matrix_0_avalon_slave_0_read,                  --                                             .read
			led_matrix_0_avalon_slave_0_readdata               => mm_interconnect_0_led_matrix_0_avalon_slave_0_readdata,              --                                             .readdata
			led_matrix_0_avalon_slave_0_writedata              => mm_interconnect_0_led_matrix_0_avalon_slave_0_writedata,             --                                             .writedata
			led_matrix_0_avalon_slave_0_byteenable             => mm_interconnect_0_led_matrix_0_avalon_slave_0_byteenable,            --                                             .byteenable
			led_matrix_0_avalon_slave_0_chipselect             => mm_interconnect_0_led_matrix_0_avalon_slave_0_chipselect,            --                                             .chipselect
			performance_checker_0_control_slave_address        => mm_interconnect_0_performance_checker_0_control_slave_address,       --          performance_checker_0_control_slave.address
			performance_checker_0_control_slave_write          => mm_interconnect_0_performance_checker_0_control_slave_write,         --                                             .write
			performance_checker_0_control_slave_readdata       => mm_interconnect_0_performance_checker_0_control_slave_readdata,      --                                             .readdata
			performance_checker_0_control_slave_writedata      => mm_interconnect_0_performance_checker_0_control_slave_writedata,     --                                             .writedata
			performance_checker_0_control_slave_begintransfer  => mm_interconnect_0_performance_checker_0_control_slave_begintransfer, --                                             .begintransfer
			pio_buttons_s1_address                             => mm_interconnect_0_pio_buttons_s1_address,                            --                               pio_buttons_s1.address
			pio_buttons_s1_write                               => mm_interconnect_0_pio_buttons_s1_write,                              --                                             .write
			pio_buttons_s1_readdata                            => mm_interconnect_0_pio_buttons_s1_readdata,                           --                                             .readdata
			pio_buttons_s1_writedata                           => mm_interconnect_0_pio_buttons_s1_writedata,                          --                                             .writedata
			pio_buttons_s1_chipselect                          => mm_interconnect_0_pio_buttons_s1_chipselect,                         --                                             .chipselect
			pio_leds_s1_address                                => mm_interconnect_0_pio_leds_s1_address,                               --                                  pio_leds_s1.address
			pio_leds_s1_write                                  => mm_interconnect_0_pio_leds_s1_write,                                 --                                             .write
			pio_leds_s1_readdata                               => mm_interconnect_0_pio_leds_s1_readdata,                              --                                             .readdata
			pio_leds_s1_writedata                              => mm_interconnect_0_pio_leds_s1_writedata,                             --                                             .writedata
			pio_leds_s1_chipselect                             => mm_interconnect_0_pio_leds_s1_chipselect,                            --                                             .chipselect
			pio_switches_s1_address                            => mm_interconnect_0_pio_switches_s1_address,                           --                              pio_switches_s1.address
			pio_switches_s1_write                              => mm_interconnect_0_pio_switches_s1_write,                             --                                             .write
			pio_switches_s1_readdata                           => mm_interconnect_0_pio_switches_s1_readdata,                          --                                             .readdata
			pio_switches_s1_writedata                          => mm_interconnect_0_pio_switches_s1_writedata,                         --                                             .writedata
			pio_switches_s1_chipselect                         => mm_interconnect_0_pio_switches_s1_chipselect,                        --                                             .chipselect
			Processor_Nios_jtag_debug_module_address           => mm_interconnect_0_processor_nios_jtag_debug_module_address,          --             Processor_Nios_jtag_debug_module.address
			Processor_Nios_jtag_debug_module_write             => mm_interconnect_0_processor_nios_jtag_debug_module_write,            --                                             .write
			Processor_Nios_jtag_debug_module_read              => mm_interconnect_0_processor_nios_jtag_debug_module_read,             --                                             .read
			Processor_Nios_jtag_debug_module_readdata          => mm_interconnect_0_processor_nios_jtag_debug_module_readdata,         --                                             .readdata
			Processor_Nios_jtag_debug_module_writedata         => mm_interconnect_0_processor_nios_jtag_debug_module_writedata,        --                                             .writedata
			Processor_Nios_jtag_debug_module_byteenable        => mm_interconnect_0_processor_nios_jtag_debug_module_byteenable,       --                                             .byteenable
			Processor_Nios_jtag_debug_module_waitrequest       => mm_interconnect_0_processor_nios_jtag_debug_module_waitrequest,      --                                             .waitrequest
			Processor_Nios_jtag_debug_module_debugaccess       => mm_interconnect_0_processor_nios_jtag_debug_module_debugaccess,      --                                             .debugaccess
			RAM_s1_address                                     => mm_interconnect_0_ram_s1_address,                                    --                                       RAM_s1.address
			RAM_s1_write                                       => mm_interconnect_0_ram_s1_write,                                      --                                             .write
			RAM_s1_readdata                                    => mm_interconnect_0_ram_s1_readdata,                                   --                                             .readdata
			RAM_s1_writedata                                   => mm_interconnect_0_ram_s1_writedata,                                  --                                             .writedata
			RAM_s1_byteenable                                  => mm_interconnect_0_ram_s1_byteenable,                                 --                                             .byteenable
			RAM_s1_chipselect                                  => mm_interconnect_0_ram_s1_chipselect,                                 --                                             .chipselect
			RAM_s1_clken                                       => mm_interconnect_0_ram_s1_clken,                                      --                                             .clken
			sysid_qsys_0_control_slave_address                 => mm_interconnect_0_sysid_qsys_0_control_slave_address,                --                   sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,               --                                             .readdata
			timer_0_s1_address                                 => mm_interconnect_0_timer_0_s1_address,                                --                                   timer_0_s1.address
			timer_0_s1_write                                   => mm_interconnect_0_timer_0_s1_write,                                  --                                             .write
			timer_0_s1_readdata                                => mm_interconnect_0_timer_0_s1_readdata,                               --                                             .readdata
			timer_0_s1_writedata                               => mm_interconnect_0_timer_0_s1_writedata,                              --                                             .writedata
			timer_0_s1_chipselect                              => mm_interconnect_0_timer_0_s1_chipselect                              --                                             .chipselect
		);

	irq_mapper : component eindopdracht_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => processor_nios_d_irq_irq        --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => processor_nios_jtag_debug_module_reset_reset, -- reset_in0.reset
			clk            => clk_clk,                                      --       clk.clk
			reset_out      => rst_controller_reset_out_reset,               -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,           --          .reset_req
			reset_req_in0  => '0',                                          -- (terminated)
			reset_in1      => '0',                                          -- (terminated)
			reset_req_in1  => '0',                                          -- (terminated)
			reset_in2      => '0',                                          -- (terminated)
			reset_req_in2  => '0',                                          -- (terminated)
			reset_in3      => '0',                                          -- (terminated)
			reset_req_in3  => '0',                                          -- (terminated)
			reset_in4      => '0',                                          -- (terminated)
			reset_req_in4  => '0',                                          -- (terminated)
			reset_in5      => '0',                                          -- (terminated)
			reset_req_in5  => '0',                                          -- (terminated)
			reset_in6      => '0',                                          -- (terminated)
			reset_req_in6  => '0',                                          -- (terminated)
			reset_in7      => '0',                                          -- (terminated)
			reset_req_in7  => '0',                                          -- (terminated)
			reset_in8      => '0',                                          -- (terminated)
			reset_req_in8  => '0',                                          -- (terminated)
			reset_in9      => '0',                                          -- (terminated)
			reset_req_in9  => '0',                                          -- (terminated)
			reset_in10     => '0',                                          -- (terminated)
			reset_req_in10 => '0',                                          -- (terminated)
			reset_in11     => '0',                                          -- (terminated)
			reset_req_in11 => '0',                                          -- (terminated)
			reset_in12     => '0',                                          -- (terminated)
			reset_req_in12 => '0',                                          -- (terminated)
			reset_in13     => '0',                                          -- (terminated)
			reset_req_in13 => '0',                                          -- (terminated)
			reset_in14     => '0',                                          -- (terminated)
			reset_req_in14 => '0',                                          -- (terminated)
			reset_in15     => '0',                                          -- (terminated)
			reset_req_in15 => '0'                                           -- (terminated)
		);

	mm_interconnect_0_jtag_debug_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_debug_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_debug_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_debug_avalon_jtag_slave_write;

	mm_interconnect_0_pio_buttons_s1_write_ports_inv <= not mm_interconnect_0_pio_buttons_s1_write;

	mm_interconnect_0_pio_switches_s1_write_ports_inv <= not mm_interconnect_0_pio_switches_s1_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_pio_leds_s1_write_ports_inv <= not mm_interconnect_0_pio_leds_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of eindopdracht
