LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY bst_7_segment IS
	PORT ( CLOCK_50 : IN STD_LOGIC;
	KEY : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
	HEX0 : OUT STD_LOGIC_VECTOR(0 TO 6);
	HEX1 : OUT STD_LOGIC_VECTOR(0 TO 6);
	HEX2 : OUT STD_LOGIC_VECTOR(0 TO 6);
	HEX3 : OUT STD_LOGIC_VECTOR(0 TO 6));
	END bst_7_segment;

ARCHITECTURE Structure OF bst_7_segment IS
	SIGNAL to_HEX : STD_LOGIC_VECTOR(31 DOWNTO 0);
	COMPONENT embedded_system IS
	PORT ( 
		clk_clk : IN STD_LOGIC;
		reset_reset_n : IN STD_LOGIC;
		to_hex_readdata: OUT STD_LOGIC_VECTOR (31 DOWNTO 0) );
	END COMPONENT embedded_system;
	
--	COMPONENT hex7seg IS
--	PORT ( hex : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
--		display : OUT STD_LOGIC_VECTOR(0 TO 6) );
--	END COMPONENT hex7seg;
BEGIN

	U0: embedded_system PORT MAP (
	clk_clk => CLOCK_50,
	reset_reset_n => KEY(0),
	to_hex_readdata(6 downto 0) => HEX0,
	to_hex_readdata(13 downto 7) => HEX1,
	to_hex_readdata(20 downto 14) => HEX2,
	to_hex_readdata(27 downto 21) => HEX3);
	
END Structure;