library ieee;
use ieee.std_logic_1164.all;

entity fsm_display is
	port (
        clk, rst: in std_ulogic;
        input1, input2, ...: in std_ulogic;
        output1, output2, ...: out std_ulogic
    );
end fsm_display;

architecture behavior of fsm_display is
   type state_type is (IDLE, SHIFT, LATCH, DISPLAY, NEXT_ROW);
	signal pr_state, nx_state: state_type;
begin

    process(clk, rst)
    begin
        if rst then
            pr_state <= idle;
        elsif rising_edge(clk) then
            pr_state <= nx_state;
        end if;
    end process;

    process(pr_state, input1, input2, ...)
    begin
        case pr_state is
          when IDLE =>
              if input1 then
                nx_state <= state1;
              else
                nx_state <= state2;
              end if;
            when SHIFT =>
                nx_state <= state2;
            when LATCH =>
                ...;
            when DISPLAY =>
                ...;
				when NEXT_ROW =>
					 ...;
        end case;
    end process;

    process(pr_state)
    begin
        case pr_state is
            when idle =>
                output1 <= '0';
                output2 <= '0';
                ... 
            when state1 =>
                output1 <= '0';
                output2 <= '1';
                ... 
            when state2 =>
                ...;
            when ... =>
                ...;
        end case;
    end process;

end architecture;